** Profile: "SCHEMATIC1-CV"  [ D:\ae\ass-SCHEMATIC1-CV.sim ] 

** Creating circuit file "ass-SCHEMATIC1-CV.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 40ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\ass-SCHEMATIC1.net" 


.END
