** Profile: "SCHEMATIC1-COMMON BASE"  [ D:\ae\common base-SCHEMATIC1-COMMON BASE.sim ] 

** Creating circuit file "common base-SCHEMATIC1-COMMON BASE.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_VCC -2 30 1 
+ LIN V_VEE 0 5 1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\common base-SCHEMATIC1.net" 


.END
