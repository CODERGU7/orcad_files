** Profile: "SCHEMATIC1-AD"  [ D:\ae\bjt-SCHEMATIC1-AD.sim ] 

** Creating circuit file "bjt-SCHEMATIC1-AD.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_VCC 0 30 1 
+ LIN V_VBB 0 5 1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\bjt-SCHEMATIC1.net" 


.END
