** Profile: "SCHEMATIC1-exp_rseries"  [ D:\ae\exp_rseries-schematic1-exp_rseries.sim ] 

** Creating circuit file "exp_rseries-schematic1-exp_rseries.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0 5 0.1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\exp_rseries-SCHEMATIC1.net" 


.END
