** Profile: "SCHEMATIC1-input"  [ D:\ae\common base-SCHEMATIC1-input.sim ] 

** Creating circuit file "common base-SCHEMATIC1-input.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_VEE 0 5 .5 
+ LIN V_VCC 0 15 5 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\common base-SCHEMATIC1.net" 


.END
