** Profile: "SCHEMATIC1-MESH"  [ D:\ae\eadtest-schematic1-mesh.sim ] 

** Creating circuit file "eadtest-schematic1-mesh.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\eadtest-SCHEMATIC1.net" 


.END
