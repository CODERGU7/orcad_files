** Profile: "SCHEMATIC1-ERA"  [ D:\ae\eadtest2-schematic1-era.sim ] 

** Creating circuit file "eadtest2-schematic1-era.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\eadtest2-SCHEMATIC1.net" 


.END
