** Profile: "SCHEMATIC1-h"  [ D:\ae\d-schematic1-h.sim ] 

** Creating circuit file "d-schematic1-h.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0 10 0.1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\d-SCHEMATIC1.net" 


.END
